// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_UART16550_CSRS_DATA_W 32
// Core Configuration Macros.
`define IOB_UART16550_CSRS_RBR_THR_DLL_ADDR 0
`define IOB_UART16550_CSRS_RBR_THR_DLL_W 8
`define IOB_UART16550_CSRS_IER_DLM_ADDR 1
`define IOB_UART16550_CSRS_IER_DLM_W 8
`define IOB_UART16550_CSRS_IIR_FCR_ADDR 2
`define IOB_UART16550_CSRS_IIR_FCR_W 8
`define IOB_UART16550_CSRS_LCR_ADDR 3
`define IOB_UART16550_CSRS_LCR_W 8
`define IOB_UART16550_CSRS_MCR_ADDR 4
`define IOB_UART16550_CSRS_MCR_W 8
`define IOB_UART16550_CSRS_LSR_ADDR 5
`define IOB_UART16550_CSRS_LSR_W 8
`define IOB_UART16550_CSRS_MSR_ADDR 6
`define IOB_UART16550_CSRS_MSR_W 8
`define IOB_UART16550_CSRS_VERSION_ADDR 8
`define IOB_UART16550_CSRS_VERSION_W 32
`define IOB_UART16550_CSRS_VERSION 24'h000104
// Core Derived Parameters. DO NOT CHANGE
`define IOB_UART16550_CSRS_ADDR_W 4
