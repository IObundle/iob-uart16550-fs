// general_operation: General operation group
// Core Constants. DO NOT CHANGE
`define TB_PBUS_SPLIT_VERSION 16'h0081
