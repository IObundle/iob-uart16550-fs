// SPDX-FileCopyrightText: 2025 IObundle
//
// SPDX-License-Identifier: MIT

`include "iob_uart16550_conf.vh"
`define IOB_CSRS_ADDR_W (`IOB_UART16550_ADDR_W+1)

