// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_UNIVERSAL_CONVERTER_IOB_WB_ADDR_W 1
`define IOB_UNIVERSAL_CONVERTER_IOB_WB_DATA_W 32
`define IOB_UNIVERSAL_CONVERTER_IOB_WB_READ_BYTES 4
// Core Configuration Macros.
`define IOB_UNIVERSAL_CONVERTER_IOB_WB_VERSION 24'h008100
