// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_UART16550_ADDR_W 5
`define IOB_UART16550_DATA_W 32
// Core Configuration Macros.
`define IOB_UART16550_VERSION 24'h000104
