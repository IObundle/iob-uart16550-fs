// general_operation: General operation group
// Core Configuration Macros.
`define IOB_LINUX_DEVICE_DRIVERS_VERSION 24'h008100
