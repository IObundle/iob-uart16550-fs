// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_IOB2WISHBONE_DATA_W 32
`define IOB_IOB2WISHBONE_ADDR_W 32
`define IOB_IOB2WISHBONE_READ_BYTES 4
// Core Configuration Macros.
`define IOB_IOB2WISHBONE_VERSION 24'h008100
