// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_UUT_ADDR_W 6
`define IOB_UUT_DATA_W 32
// Core Configuration Macros.
`define IOB_UUT_VERSION 24'h008100
