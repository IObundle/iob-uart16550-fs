// general_operation: General operation group
// Core Configuration Macros.
`define IOB_UART16550_ST_VERSION 24'h008100
